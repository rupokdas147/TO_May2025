* Extracted by KLayout with SG13G2 LVS runset on : 09/05/2025 17:10

.SUBCKT FMD_QNC_60_GHZ_LA
C$1 \$I328611 \$1 cap_cmim w=30u l=30u A=900p P=120u m=16
C$9 \$I328612 \$1 cap_cmim w=30u l=30u A=900p P=120u m=6
C$21 \$I328629 \$1 cap_cmim w=30u l=30u A=900p P=120u m=2
C$23 \$I328637 \$1 cap_cmim w=30u l=30u A=900p P=120u m=2
C$25 \$I328638 \$1 cap_cmim w=30u l=30u A=900p P=120u m=2
C$29 \$I328648 \$1 cap_cmim w=30u l=30u A=900p P=120u m=2
R$31 \$I328629 \$I328631 rsil w=20u l=22u ps=0 b=0 m=1
R$32 \$I328629 \$I328630 rsil w=20u l=22u ps=0 b=0 m=1
R$33 \$I328613 \$I328611 rppd w=18u l=2.7u ps=0 b=0 m=1
R$34 \$I328614 \$I328611 rppd w=18u l=2.7u ps=0 b=0 m=1
R$35 \$I328639 \$1 rsil w=20u l=18u ps=0 b=0 m=2
R$37 \$I328618 \$I328634 rppd w=18u l=2u ps=0 b=0 m=1
R$38 \$I328617 \$I328643 rppd w=18u l=2u ps=0 b=0 m=1
R$39 \$I328633 \$1 rsil w=20u l=2.6u ps=0 b=0 m=2
R$41 \$1 \$I328641 rsil w=20u l=2.6u ps=0 b=0 m=2
R$43 \$I328634 \$I328611 rppd w=21u l=2u ps=0 b=0 m=1
R$44 \$I328643 \$I328611 rppd w=21u l=2u ps=0 b=0 m=1
Q$45 \$I328638 \$I328612 \$I328639 \$1 npn13G2 AE=0.063p PE=1.94u AB=19.2965p
+ PB=19.32u AC=19.283334p PC=19.31u NE=3 m=3
R$48 \$I328636 \$I328635 rppd w=12u l=3.1u ps=0 b=0 m=1
R$49 \$I328640 \$I328642 rppd w=12u l=3.1u ps=0 b=0 m=1
R$50 \$I328644 \$I328611 rppd w=5u l=13u ps=0 b=0 m=1
C$51 \$I328647 \$1 cap_cmim w=30u l=30u A=900p P=120u m=1
R$52 \$I328615 \$I328647 rsil w=2u l=10.38u ps=0 b=0 m=1
R$53 \$I328616 \$I328647 rsil w=2u l=10.38u ps=0 b=0 m=1
R$54 \$1 \$I328649 rsil w=20u l=3.2u ps=0 b=0 m=2
R$56 \$I328648 \$I328619 rppd w=12u l=3.3u ps=0 b=0 m=1
R$57 \$I328648 \$I328620 rppd w=12u l=3.3u ps=0 b=0 m=1
Q$58 \$I328632 \$I328612 \$I328633 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q$68 \$I328629 \$I328629 \$I328632 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q$78 \$I328637 \$I328612 \$I328641 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q$88 \$I328611 \$I328611 \$I328646 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q$98 \$I328648 \$I328612 \$I328649 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q$108 \$I328611 \$I328611 \$I328650 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q$118 \$I328614 \$I328618 \$I328631 \$1 npn13G2 AE=0.063p PE=1.94u AB=31.9135p
+ PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
Q$123 \$I328613 \$I328617 \$I328630 \$1 npn13G2 AE=0.063p PE=1.94u AB=31.9135p
+ PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
Q$128 \$I328617 \$I328640 \$I328637 \$1 npn13G2 AE=0.063p PE=1.94u AB=31.9135p
+ PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
Q$133 \$I328618 \$I328636 \$I328637 \$1 npn13G2 AE=0.063p PE=1.94u AB=31.9135p
+ PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
Q$138 \$I328646 \$I328616 \$I328620 \$1 npn13G2 AE=0.063p PE=1.94u AB=31.9135p
+ PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
Q$143 \$I328650 \$I328615 \$I328619 \$1 npn13G2 AE=0.063p PE=1.94u AB=31.9135p
+ PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
R$148 \$I328647 \$I328611 rhigh w=2u l=4u ps=0 b=0 m=2
R$150 \$I328654 \$I328647 rhigh w=4u l=4u ps=0 b=0 m=1
R$151 \$I328652 \$I328653 rhigh w=4u l=4u ps=0 b=0 m=1
R$152 \$I328655 \$I328652 rhigh w=2u l=6.4u ps=0 b=0 m=2
Q$154 \$I328636 \$I328620 \$I328638 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
Q$155 \$I328611 \$I328643 \$I328642 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
Q$156 \$I328640 \$I328619 \$I328638 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
Q$157 \$I328611 \$I328634 \$I328635 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
Q$158 \$I328645 \$I328644 \$I328612 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
Q$159 \$I328644 \$I328612 \$1 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
Q$160 \$I328611 \$I328611 \$I328645 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
Q$161 \$I328647 \$I328654 \$I328655 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
Q$162 \$I328652 \$I328653 \$1 \$1 npn13G2 AE=0.063p PE=1.94u AB=6.6795p
+ PB=11.92u AC=6.670034p PC=11.91u NE=1 m=1
.ENDS FMD_QNC_60_GHZ_LA
